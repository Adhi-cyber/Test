module buffer_gate(
	input d,
	input e,
	output y);

and(y,d,e);

endmodule
