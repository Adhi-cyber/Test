module and_gate_des(
	input a,
	input b,
	output c);

and(c,a,b);

endmodule
