module and_gate_ass(
	input a,
	input b,
	output c);

assign c = a&b;
endmodule
